interface dut_if;

logic        clk;
logic [31:0] addr;
logic [31:0] data;
logic [31:0] delay;

endinterface