`define TIMEOUT 1000000
