//------------------------------------------------------------
//   Copyright 2010-2011 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

module mem_ss_wrapper(interface AHB);

mem_ss u_1(.HCLK(AHB.HCLK),
           .HRESETn(AHB.HRESETn),
           .HADDR(AHB.HADDR[30:0]),
           .HWRITE(AHB.HWRITE),
           .HTRANS(AHB.HTRANS),
           .HSIZE(AHB.HSIZE),
           .HBURST(AHB.HBURST),
           .HPROT(AHB.HPROT),
           .HWDATA(AHB.HWDATA),
           .HSEL(AHB.HSEL),
           .HREADY(AHB.HREADY),
           .HRDATA(AHB.HRDATA),
           .HRESP(AHB.HRESP)
             );

endmodule: mem_ss_wrapper