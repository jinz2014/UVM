../ipxact/uart_ctrl_regs.sv